module audio_main (
	CLOCK_50,
	KEY,
	AUD_ADCDAT,

	AUD_BCLK,
	AUD_ADCLRCK,
	AUD_DACLRCK,

	FPGA_I2C_SDAT,

	AUD_XCK,
	AUD_DACDAT,

	FPGA_I2C_SCLK,
	SW,
);

input				CLOCK_50;
input		[3:0]	KEY;
input		[3:0]	SW;
reg [1:0] sound_sel;

input				AUD_ADCDAT;

inout				AUD_BCLK;
inout				AUD_ADCLRCK;
inout				AUD_DACLRCK;
inout				FPGA_I2C_SDAT;
output				AUD_XCK;
output				AUD_DACDAT;
output				FPGA_I2C_SCLK;


wire				audio_in_available;
wire		[31:0]	left_channel_audio_in;
wire		[31:0]	right_channel_audio_in;
wire				read_audio_in;
wire [5:0]	audio_from_ram;
wire				audio_out_allowed;
wire		[31:0]	left_channel_audio_out;
wire		[31:0]	right_channel_audio_out;
wire				write_audio_out;
wire [17:0] address_count;

reg [18:0] delay_cnt;
wire [18:0] delay;
reg [13:0] addr_count, soundstart, soundend;;
reg [10:0] clock_count;
reg snd;


reg [22:0] beatCountMario;
reg [9:0] addressMario; 
													
sound_rom r1(.address(addressMario), .clock(CLOCK_50), .q(delay));
win_rom w1(.address(addressMario), .clock(CLOCK_50), .q(delay));

always @(*) begin
    if (~SW[0]) begin
        sound_sel <= 2'b00; // Mario sound
    end else if (~SW[1]) begin
        sound_sel <= 2'b01; // Win sound
    end else begin
        sound_sel <= 2'b10; // Default or other sound
    end
end

always @(posedge CLOCK_50)
	if(delay_cnt == delay) begin
		delay_cnt <= 0;
		snd <= !snd;
	end else delay_cnt <= delay_cnt + 1;


always @(posedge CLOCK_50) begin
	case(sound_sel)
		2'b00: begin //mario sound 
		if(beatCountMario == 23'd2500000)begin
			beatCountMario <= 23'b0;
			if(addressMario < 10'd999)
				addressMario <= addressMario + 1;
			else begin
				addressMario <= 0;
				beatCountMario <= 0;
			end
		end
		else 
			beatCountMario <= beatCountMario + 1;
		end

		2'b01: begin //win sound 
			soundstart <= 18'd0; //
			soundend <= 18'd16395;

			if (clock_count == 11'd1200) begin
				if (addr_count == soundend) begin 
					addr_count <= soundstart;
				end
				else if ((addr_count >= soundstart) && (addr_count < soundend)) begin
					addr_count <= addr_count + 1'b1;
					clock_count <= 0;
				end
				else addr_count <= soundstart;
			end
		else clock_count <= clock_count + 1;
		end

		default: begin
		end
	endcase
end

wire [31:0] sound = snd ? 32'd100000000 : -32'd100000000;
assign address_count = addr_count;

assign read_audio_in			= audio_in_available & audio_out_allowed;
assign left_channel_audio_out	= left_channel_audio_in+sound;
assign right_channel_audio_out	= left_channel_audio_in+sound;
assign write_audio_out			= audio_in_available & audio_out_allowed;

Audio_Controller Audio_Controller (
	.CLOCK_50					(CLOCK_50),
	.reset						(~KEY[0]),
	.clear_audio_in_memory	(),
	.read_audio_in				(read_audio_in),
	.clear_audio_out_memory		(),
	.left_channel_audio_out		(left_channel_audio_out),
	.right_channel_audio_out	(right_channel_audio_out),
	.write_audio_out			(1'b1),
	.AUD_ADCDAT					(AUD_ADCDAT),
	.AUD_BCLK					(AUD_BCLK),
	.AUD_ADCLRCK				(AUD_ADCLRCK),
	.AUD_DACLRCK				(AUD_DACLRCK),
	.audio_in_available			(audio_in_available),
	.left_channel_audio_in		(left_channel_audio_in),
	.right_channel_audio_in		(right_channel_audio_in),
	.audio_out_allowed			(audio_out_allowed),
	.AUD_XCK					(AUD_XCK),
	.AUD_DACDAT					(AUD_DACDAT)

);

avconf #(.USE_MIC_INPUT(1)) avc (
	.FPGA_I2C_SCLK					(FPGA_I2C_SCLK),
	.FPGA_I2C_SDAT					(FPGA_I2C_SDAT),
	.CLOCK_50					(CLOCK_50),
	.reset						(~KEY[0])
);
endmodule