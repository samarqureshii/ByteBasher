module final() //ful system integration

fill annie();
endmodule