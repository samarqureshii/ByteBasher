module final() //system level integration 
endmodule