module moduleName (
    ports
);
endmodule